module fantasticfft_top #(
    parameter NUM_POINTS = 8
) (
    input logic clk
);
    
endmodule