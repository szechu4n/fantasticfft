`timescale 1 ns/100 ps

`include "rtl/fixedpoint.sv"

module sine_lut (
   input  logic [5 : 0] start,
   input  logic [5 : 0] step,
   output logic signed [15 : 0] out [0 : 7]
);

always_comb begin : lut
   int i;
   for (i = 0; i < 8; i = i + 1) begin
      case (start + i * step)
         6'h00: out[i] = $sin(2 * 3.1415926 * 0  / 64) * 2**8;
         6'h01: out[i] = $sin(2 * 3.1415926 * 1  / 64) * 2**8; 
         6'h02: out[i] = $sin(2 * 3.1415926 * 2  / 64) * 2**8;
         6'h03: out[i] = $sin(2 * 3.1415926 * 3  / 64) * 2**8;
         6'h04: out[i] = $sin(2 * 3.1415926 * 4  / 64) * 2**8;
         6'h05: out[i] = $sin(2 * 3.1415926 * 5  / 64) * 2**8;
         6'h06: out[i] = $sin(2 * 3.1415926 * 6  / 64) * 2**8;
         6'h07: out[i] = $sin(2 * 3.1415926 * 7  / 64) * 2**8;
         6'h08: out[i] = $sin(2 * 3.1415926 * 8  / 64) * 2**8;
         6'h09: out[i] = $sin(2 * 3.1415926 * 9  / 64) * 2**8;
         6'h0a: out[i] = $sin(2 * 3.1415926 * 10 / 64) * 2**8;
         6'h0b: out[i] = $sin(2 * 3.1415926 * 11 / 64) * 2**8;
         6'h0c: out[i] = $sin(2 * 3.1415926 * 12 / 64) * 2**8;
         6'h0d: out[i] = $sin(2 * 3.1415926 * 13 / 64) * 2**8;
         6'h0e: out[i] = $sin(2 * 3.1415926 * 14 / 64) * 2**8;
         6'h0f: out[i] = $sin(2 * 3.1415926 * 15 / 64) * 2**8;
         6'h10: out[i] = $sin(2 * 3.1415926 * 16 / 64) * 2**8;
         6'h11: out[i] = $sin(2 * 3.1415926 * 17 / 64) * 2**8;
         6'h12: out[i] = $sin(2 * 3.1415926 * 18 / 64) * 2**8;
         6'h13: out[i] = $sin(2 * 3.1415926 * 19 / 64) * 2**8;
         6'h14: out[i] = $sin(2 * 3.1415926 * 20 / 64) * 2**8;
         6'h15: out[i] = $sin(2 * 3.1415926 * 21 / 64) * 2**8;
         6'h16: out[i] = $sin(2 * 3.1415926 * 22 / 64) * 2**8;
         6'h17: out[i] = $sin(2 * 3.1415926 * 23 / 64) * 2**8;
         6'h18: out[i] = $sin(2 * 3.1415926 * 24 / 64) * 2**8;
         6'h19: out[i] = $sin(2 * 3.1415926 * 25 / 64) * 2**8;
         6'h1a: out[i] = $sin(2 * 3.1415926 * 26 / 64) * 2**8;
         6'h1b: out[i] = $sin(2 * 3.1415926 * 27 / 64) * 2**8;
         6'h1c: out[i] = $sin(2 * 3.1415926 * 28 / 64) * 2**8;
         6'h1d: out[i] = $sin(2 * 3.1415926 * 29 / 64) * 2**8;
         6'h1e: out[i] = $sin(2 * 3.1415926 * 30 / 64) * 2**8;
         6'h1f: out[i] = $sin(2 * 3.1415926 * 31 / 64) * 2**8;
         6'h20: out[i] = $sin(2 * 3.1415926 * 32 / 64) * 2**8;
         6'h21: out[i] = $sin(2 * 3.1415926 * 33 / 64) * 2**8;
         6'h22: out[i] = $sin(2 * 3.1415926 * 34 / 64) * 2**8;
         6'h23: out[i] = $sin(2 * 3.1415926 * 35 / 64) * 2**8;
         6'h24: out[i] = $sin(2 * 3.1415926 * 36 / 64) * 2**8;
         6'h25: out[i] = $sin(2 * 3.1415926 * 37 / 64) * 2**8;
         6'h26: out[i] = $sin(2 * 3.1415926 * 38 / 64) * 2**8;
         6'h27: out[i] = $sin(2 * 3.1415926 * 39 / 64) * 2**8;
         6'h28: out[i] = $sin(2 * 3.1415926 * 40 / 64) * 2**8;
         6'h29: out[i] = $sin(2 * 3.1415926 * 41 / 64) * 2**8;
         6'h2a: out[i] = $sin(2 * 3.1415926 * 42 / 64) * 2**8;
         6'h2b: out[i] = $sin(2 * 3.1415926 * 43 / 64) * 2**8;
         6'h2c: out[i] = $sin(2 * 3.1415926 * 44 / 64) * 2**8;
         6'h2d: out[i] = $sin(2 * 3.1415926 * 45 / 64) * 2**8;
         6'h2e: out[i] = $sin(2 * 3.1415926 * 46 / 64) * 2**8;
         6'h2f: out[i] = $sin(2 * 3.1415926 * 47 / 64) * 2**8;
         6'h30: out[i] = $sin(2 * 3.1415926 * 48 / 64) * 2**8;
         6'h31: out[i] = $sin(2 * 3.1415926 * 49 / 64) * 2**8;
         6'h32: out[i] = $sin(2 * 3.1415926 * 50 / 64) * 2**8;
         6'h33: out[i] = $sin(2 * 3.1415926 * 51 / 64) * 2**8;
         6'h34: out[i] = $sin(2 * 3.1415926 * 52 / 64) * 2**8;
         6'h35: out[i] = $sin(2 * 3.1415926 * 53 / 64) * 2**8;
         6'h36: out[i] = $sin(2 * 3.1415926 * 54 / 64) * 2**8;
         6'h37: out[i] = $sin(2 * 3.1415926 * 55 / 64) * 2**8;
         6'h38: out[i] = $sin(2 * 3.1415926 * 56 / 64) * 2**8;
         6'h39: out[i] = $sin(2 * 3.1415926 * 57 / 64) * 2**8;
         6'h3a: out[i] = $sin(2 * 3.1415926 * 58 / 64) * 2**8;
         6'h3b: out[i] = $sin(2 * 3.1415926 * 59 / 64) * 2**8;
         6'h3c: out[i] = $sin(2 * 3.1415926 * 60 / 64) * 2**8;
         6'h3d: out[i] = $sin(2 * 3.1415926 * 61 / 64) * 2**8;
         6'h3e: out[i] = $sin(2 * 3.1415926 * 62 / 64) * 2**8;
         6'h3f: out[i] = $sin(2 * 3.1415926 * 63 / 64) * 2**8;
      endcase
   end
end

endmodule

module cosine_lut (
   input  logic [5 : 0] start,
   input  logic [5 : 0] step,
   output logic signed [15 : 0] out [0 : 7]
);

always_comb begin : lut
   int i;
   for (i = 0; i < 8; i = i + 1) begin
      case (start + i * step)
         6'h00: out[i] = $cos(2 * 3.1415926 * 0  / 64) * 2**8;
         6'h01: out[i] = $cos(2 * 3.1415926 * 1  / 64) * 2**8; 
         6'h02: out[i] = $cos(2 * 3.1415926 * 2  / 64) * 2**8;
         6'h03: out[i] = $cos(2 * 3.1415926 * 3  / 64) * 2**8;
         6'h04: out[i] = $cos(2 * 3.1415926 * 4  / 64) * 2**8;
         6'h05: out[i] = $cos(2 * 3.1415926 * 5  / 64) * 2**8;
         6'h06: out[i] = $cos(2 * 3.1415926 * 6  / 64) * 2**8;
         6'h07: out[i] = $cos(2 * 3.1415926 * 7  / 64) * 2**8;
         6'h08: out[i] = $cos(2 * 3.1415926 * 8  / 64) * 2**8;
         6'h09: out[i] = $cos(2 * 3.1415926 * 9  / 64) * 2**8;
         6'h0a: out[i] = $cos(2 * 3.1415926 * 10 / 64) * 2**8;
         6'h0b: out[i] = $cos(2 * 3.1415926 * 11 / 64) * 2**8;
         6'h0c: out[i] = $cos(2 * 3.1415926 * 12 / 64) * 2**8;
         6'h0d: out[i] = $cos(2 * 3.1415926 * 13 / 64) * 2**8;
         6'h0e: out[i] = $cos(2 * 3.1415926 * 14 / 64) * 2**8;
         6'h0f: out[i] = $cos(2 * 3.1415926 * 15 / 64) * 2**8;
         6'h10: out[i] = $cos(2 * 3.1415926 * 16 / 64) * 2**8;
         6'h11: out[i] = $cos(2 * 3.1415926 * 17 / 64) * 2**8;
         6'h12: out[i] = $cos(2 * 3.1415926 * 18 / 64) * 2**8;
         6'h13: out[i] = $cos(2 * 3.1415926 * 19 / 64) * 2**8;
         6'h14: out[i] = $cos(2 * 3.1415926 * 20 / 64) * 2**8;
         6'h15: out[i] = $cos(2 * 3.1415926 * 21 / 64) * 2**8;
         6'h16: out[i] = $cos(2 * 3.1415926 * 22 / 64) * 2**8;
         6'h17: out[i] = $cos(2 * 3.1415926 * 23 / 64) * 2**8;
         6'h18: out[i] = $cos(2 * 3.1415926 * 24 / 64) * 2**8;
         6'h19: out[i] = $cos(2 * 3.1415926 * 25 / 64) * 2**8;
         6'h1a: out[i] = $cos(2 * 3.1415926 * 26 / 64) * 2**8;
         6'h1b: out[i] = $cos(2 * 3.1415926 * 27 / 64) * 2**8;
         6'h1c: out[i] = $cos(2 * 3.1415926 * 28 / 64) * 2**8;
         6'h1d: out[i] = $cos(2 * 3.1415926 * 29 / 64) * 2**8;
         6'h1e: out[i] = $cos(2 * 3.1415926 * 30 / 64) * 2**8;
         6'h1f: out[i] = $cos(2 * 3.1415926 * 31 / 64) * 2**8;
         6'h20: out[i] = $cos(2 * 3.1415926 * 32 / 64) * 2**8;
         6'h21: out[i] = $cos(2 * 3.1415926 * 33 / 64) * 2**8;
         6'h22: out[i] = $cos(2 * 3.1415926 * 34 / 64) * 2**8;
         6'h23: out[i] = $cos(2 * 3.1415926 * 35 / 64) * 2**8;
         6'h24: out[i] = $cos(2 * 3.1415926 * 36 / 64) * 2**8;
         6'h25: out[i] = $cos(2 * 3.1415926 * 37 / 64) * 2**8;
         6'h26: out[i] = $cos(2 * 3.1415926 * 38 / 64) * 2**8;
         6'h27: out[i] = $cos(2 * 3.1415926 * 39 / 64) * 2**8;
         6'h28: out[i] = $cos(2 * 3.1415926 * 40 / 64) * 2**8;
         6'h29: out[i] = $cos(2 * 3.1415926 * 41 / 64) * 2**8;
         6'h2a: out[i] = $cos(2 * 3.1415926 * 42 / 64) * 2**8;
         6'h2b: out[i] = $cos(2 * 3.1415926 * 43 / 64) * 2**8;
         6'h2c: out[i] = $cos(2 * 3.1415926 * 44 / 64) * 2**8;
         6'h2d: out[i] = $cos(2 * 3.1415926 * 45 / 64) * 2**8;
         6'h2e: out[i] = $cos(2 * 3.1415926 * 46 / 64) * 2**8;
         6'h2f: out[i] = $cos(2 * 3.1415926 * 47 / 64) * 2**8;
         6'h30: out[i] = $cos(2 * 3.1415926 * 48 / 64) * 2**8;
         6'h31: out[i] = $cos(2 * 3.1415926 * 49 / 64) * 2**8;
         6'h32: out[i] = $cos(2 * 3.1415926 * 50 / 64) * 2**8;
         6'h33: out[i] = $cos(2 * 3.1415926 * 51 / 64) * 2**8;
         6'h34: out[i] = $cos(2 * 3.1415926 * 52 / 64) * 2**8;
         6'h35: out[i] = $cos(2 * 3.1415926 * 53 / 64) * 2**8;
         6'h36: out[i] = $cos(2 * 3.1415926 * 54 / 64) * 2**8;
         6'h37: out[i] = $cos(2 * 3.1415926 * 55 / 64) * 2**8;
         6'h38: out[i] = $cos(2 * 3.1415926 * 56 / 64) * 2**8;
         6'h39: out[i] = $cos(2 * 3.1415926 * 57 / 64) * 2**8;
         6'h3a: out[i] = $cos(2 * 3.1415926 * 58 / 64) * 2**8;
         6'h3b: out[i] = $cos(2 * 3.1415926 * 59 / 64) * 2**8;
         6'h3c: out[i] = $cos(2 * 3.1415926 * 60 / 64) * 2**8;
         6'h3d: out[i] = $cos(2 * 3.1415926 * 61 / 64) * 2**8;
         6'h3e: out[i] = $cos(2 * 3.1415926 * 62 / 64) * 2**8;
         6'h3f: out[i] = $cos(2 * 3.1415926 * 63 / 64) * 2**8;
      endcase
   end
end

endmodule