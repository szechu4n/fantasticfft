module fantasticfft_ram #(
    parameter DEPTH = 64
) (
    input logic clk,
    input logic reset,
    input logic addr_a,
    input logic addr_b,
    input logic wr_a,
    input logic wr_b
    
);
    
endmodule