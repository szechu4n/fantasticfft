`timescale 1ns/10ps

// Andrew Sweeney
// CPE 527 Lab 004
// Multiplier Test Bench

// verilator lint_off all


module fantastic_fft8_tb (
    fantasticfft_fft8_if fft8if
);
    initial begin
        $finish();
    end
endmodule
